`timescale 1ns/1ps
//15 MHz Clock / 115200 = 130 baud rate
module top();
	parameter clocks_per_bit = 130;

	reg clk = 0;
	reg t_data_valid = 0;
	wire t_active;
	wire u_operation;
	reg [7:0] t_parallel_data = 0;
	wire t_serial_data;
	wire [7:0] r_parallel_data;
	wire r_data_valid;
	wire t_complete;

	u_receiver #(.clocks_per_bit(clocks_per_bit)) 
		uri (.clk(clk), .serial_data(u_operation), .data_valid(r_data_valid), .parallel_data(r_parallel_data));
	
	u_transmitter #(.clocks_per_bit(clocks_per_bit))
		uti (.clk(clk), .parallel_data(t_parallel_data), .data_valid(t_data_valid), .active(t_active), .serial_data(t_serial_data), .complete(t_complete));

	assign u_operation = t_active ? t_serial_data : 1'b1; //when the transmitter is not active, uart recieve operation is high
	
	always 
		#20 clk <= !clk;
	
	initial begin
		@(posedge clk);
		t_data_valid = 1'b1;
		t_parallel_data = 8'd37;
		@(posedge clk);
		t_data_valid = 1'b0;
		
		@(posedge r_data_valid);
		if(r_parallel_data == 8'd37)
			$display("Correct data");
		else
			$display("Incorrect data");
		$finish();
	end
endmodule
			